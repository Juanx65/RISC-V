// Project timescale
`timescale 1ns / 1ps